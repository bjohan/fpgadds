library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

entity lookup_table is
    	port ( 
		clk : in  STD_LOGIC;
	
		x 	: in std_logic_vector(6 - 1 downto 0);
		y	: out std_logic_vector(12 - 1 downto 0)
           	);
end lookup_table;

architecture Behavioral of lookup_table is
begin
	p_coount : process(clk)
	begin
		if rising_edge(clk) then

			case x is
				when "000000" => y <= "000000000000";
				when "000001" => y <= "000001100110";
				when "000010" => y <= "000011001100";
				when "000011" => y <= "000100110010";
				when "000100" => y <= "000110010111";
				when "000101" => y <= "000111111101";
				when "000110" => y <= "001001100010";
				when "000111" => y <= "001011000111";
				when "001000" => y <= "001100101011";
				when "001001" => y <= "001110001111";
				when "001010" => y <= "001111110010";
				when "001011" => y <= "010001010101";
				when "001100" => y <= "010010110111";
				when "001101" => y <= "010100011000";
				when "001110" => y <= "010101111000";
				when "001111" => y <= "010111011000";
				when "010000" => y <= "011000110110";
				when "010001" => y <= "011010010100";
				when "010010" => y <= "011011110000";
				when "010011" => y <= "011101001100";
				when "010100" => y <= "011110100110";
				when "010101" => y <= "011111111111";
				when "010110" => y <= "100001010111";
				when "010111" => y <= "100010101101";
				when "011000" => y <= "100100000010";
				when "011001" => y <= "100101010110";
				when "011010" => y <= "100110101000";
				when "011011" => y <= "100111111001";
				when "011100" => y <= "101001001000";
				when "011101" => y <= "101010010101";
				when "011110" => y <= "101011100001";
				when "011111" => y <= "101100101011";
				when "100000" => y <= "101101110011";
				when "100001" => y <= "101110111001";
				when "100010" => y <= "101111111110";
				when "100011" => y <= "110001000000";
				when "100100" => y <= "110010000001";
				when "100101" => y <= "110011000000";
				when "100110" => y <= "110011111100";
				when "100111" => y <= "110100110111";
				when "101000" => y <= "110101101111";
				when "101001" => y <= "110110100110";
				when "101010" => y <= "110111011010";
				when "101011" => y <= "111000001100";
				when "101100" => y <= "111000111100";
				when "101101" => y <= "111001101001";
				when "101110" => y <= "111010010100";
				when "101111" => y <= "111010111101";
				when "110000" => y <= "111011100011";
				when "110001" => y <= "111100001000";
				when "110010" => y <= "111100101001";
				when "110011" => y <= "111101001001";
				when "110100" => y <= "111101100101";
				when "110101" => y <= "111110000000";
				when "110110" => y <= "111110011000";
				when "110111" => y <= "111110101101";
				when "111000" => y <= "111111000000";
				when "111001" => y <= "111111010001";
				when "111010" => y <= "111111011111";
				when "111011" => y <= "111111101010";
				when "111100" => y <= "111111110011";
				when "111101" => y <= "111111111001";
				when "111110" => y <= "111111111101";
				when "111111" => y <= "111111111111";
				when others => y <= (others => '0');

			end case;
		end if;
	end process;

end Behavioral;
