----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:40:53 08/24/2016 
-- Design Name: 
-- Module Name:    tb - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity tb is
end tb;

architecture Behavioral of tb is
component dds_papilio_pro_top_str
    Port ( clk : in  STD_LOGIC;
           led1 : out  STD_LOGIC);
end component;


signal clk  : std_logic:= '0';
signal led : std_logic;

begin
i_top : dds_papilio_pro_top_str
port map(clk => clk, led1 => led);

end Behavioral;

